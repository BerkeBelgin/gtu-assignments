module and32b(out,i1,i0);
input [31:0] i1, i0;
output [31:0] out;

and a0(out[0],i1[0],i0[0]);
and a1(out[1],i1[1],i0[1]);
and a2(out[2],i1[2],i0[2]);
and a3(out[3],i1[3],i0[3]);
and a4(out[4],i1[4],i0[4]);
and a5(out[5],i1[5],i0[5]);
and a6(out[6],i1[6],i0[6]);
and a7(out[7],i1[7],i0[7]);
and a8(out[8],i1[8],i0[8]);
and a9(out[9],i1[9],i0[9]);
and a10(out[10],i1[10],i0[10]);
and a11(out[11],i1[11],i0[11]);
and a12(out[12],i1[12],i0[12]);
and a13(out[13],i1[13],i0[13]);
and a14(out[14],i1[14],i0[14]);
and a15(out[15],i1[15],i0[15]);
and a16(out[16],i1[16],i0[16]);
and a17(out[17],i1[17],i0[17]);
and a18(out[18],i1[18],i0[18]);
and a19(out[19],i1[19],i0[19]);
and a20(out[20],i1[20],i0[20]);
and a21(out[21],i1[21],i0[21]);
and a22(out[22],i1[22],i0[22]);
and a23(out[23],i1[23],i0[23]);
and a24(out[24],i1[24],i0[24]);
and a25(out[25],i1[25],i0[25]);
and a26(out[26],i1[26],i0[26]);
and a27(out[27],i1[27],i0[27]);
and a28(out[28],i1[28],i0[28]);
and a29(out[29],i1[29],i0[29]);
and a30(out[30],i1[30],i0[30]);
and a31(out[31],i1[31],i0[31]);

endmodule
